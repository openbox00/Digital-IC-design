module lcd_ctrl(clk, reset, datain, cmd, cmd_valid, dataout, output_valid, busy);
input clk;
input reset;
input [7:0] datain;
input [2:0] cmd;
input cmd_valid;
output [7:0] dataout;
output output_valid;
output busy;
