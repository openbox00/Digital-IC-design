`timescale 1ns/10ps

module simple_alu(
        opcode,
        in1,
        in2,
        overflow,
        result
        );

input   [2:0]   opcode;    
input   [3:0]   in1;
input   [3:0]   in2;
output          overflow;
output  [3:0]   result;

/*---------------------------------------
              Your Code
---------------------------------------*/
endmodule