`timescale 1ns/10ps

module Mask(
		data_out,
		out_valid,
		busy,
		data_in,
		clk,
		rst
        );
output [7:0] data_out;
output out_valid;
output busy;
input [7:0] data_in;
input clk;
input rst;

/*---------------------------------------
              Your Code
---------------------------------------*/

endmodule
